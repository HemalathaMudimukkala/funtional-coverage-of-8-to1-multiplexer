module tb;
  reg a,b,c,d,e,f,g,h;
  reg [2:0] sel;
  wire y;
  
  mux dut(a,b,c,d,e,f,g,h,sel,y);
  
  covergroup cvr_mux;
    option.per_instance=1;
    
    coverpoint a{
      bins a_l = {0};
      bins a_h = {1};
    }
    
    coverpoint b{
      bins b_l = {0};
      bins b_h = {1};
    }
    
    coverpoint c{
      bins c_l = {0};
      bins c_h = {1};
    }
    
    coverpoint d{
      bins d_l = {0};
      bins d_h = {1};
    }
    
    coverpoint e{
      bins e_l = {0};
      bins e_h = {1};
    }
    
    coverpoint f{
      bins f_l = {0};
      bins f_h = {1};
    }
    
    coverpoint g{
      bins g_l = {0};
      bins g_h = {1};
    }
    
    coverpoint h{
      bins h_l = {0};
      bins h_h = {1};
    }
    coverpoint sel;
    coverpoint y{
      bins y_l = {0};
      bins y_h = {1};
    }
    
    cross_a_sel: cross sel,a{
      ignore_bins sel_a = binsof(sel)intersect{[1:7]};
    }
    cross_b_sel: cross sel,b{
      ignore_bins sel_b = binsof(sel)intersect{0,[2:7]};
    }
    cross_c_sel: cross sel,c{
      ignore_bins sel_c = binsof(sel)intersect{0,1,[3:7]};
    }
    cross_d_sel: cross sel,d{
      ignore_bins sel_d = binsof(sel)intersect{[0:2],[4:7]};
    }
    cross_e_sel: cross sel,e{
      ignore_bins sel_e = binsof(sel)intersect{[0:3],[5:7]};
    }
    cross_f_sel: cross sel,f{
      ignore_bins sel_f = binsof(sel)intersect{[0:4],6,7};
    }
    cross_g_sel: cross sel,g{
      ignore_bins sel_g = binsof(sel)intersect{[0:5],7};
    }
    cross_h_sel: cross sel,h{
      ignore_bins sel_h = binsof(sel)intersect{[0:6]};
    }
    
 
   endgroup
   
  cvr_mux cvm = new();
  
  initial begin
    for(int i=0;i<100; i++) begin
      sel = $urandom();
      {a,b,c,d,e,f,g,h} = $urandom();
      cvm.sample();
      #10;
    end
  end
  
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars;
    #1200;
    $finish;
  end
  
endmodule
